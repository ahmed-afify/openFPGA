//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: FPGA Verilog Testbench for Top-level netlist of Design: and2
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Tue Aug  4 14:48:13 2020
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

module and2_autocheck_top_tb;
// ----- Local wires for global ports of FPGA fabric -----
wire [0:0] pReset;
wire [0:0] prog_clk;
wire [0:0] set;
wire [0:0] reset;
wire [0:0] clk;

// ----- Local wires for I/Os of FPGA fabric -----
wire [0:63] gfpga_pad_iopad_pad;



reg [0:0] config_done;
wire [0:0] prog_clock;
reg [0:0] prog_clock_reg;
wire [0:0] op_clock;
reg [0:0] op_clock_reg;
reg [0:0] prog_reset;
reg [0:0] prog_set;
reg [0:0] greset;
reg [0:0] gset;
// ---- Configuration-chain head -----
reg [0:0] ccff_head;
// ---- Configuration-chain tail -----
wire [0:0] ccff_tail;
// ----- Shared inputs -------
	reg [0:0] a;
	reg [0:0] b;

// ----- FPGA fabric outputs -------
	wire [0:0] out_c_fpga;

`ifdef AUTOCHECKED_SIMULATION

// ----- Benchmark outputs -------
	wire [0:0] out_c_benchmark;

// ----- Output vectors checking flags -------
	reg [0:0] out_c_flag;

`endif

// ----- Error counter -----
	integer nb_error= 0;
// ----- Number of clock cycles in configuration phase: 1877 -----
// ----- Begin configuration done signal generation -----
initial
	begin
		config_done[0] = {1{1'b0}};
	end

// ----- End configuration done signal generation -----

// ----- Begin raw programming clock signal generation -----
initial
	begin
		prog_clock_reg[0] = {1{1'b0}};
	end
always
	begin
		#5	prog_clock_reg[0] = ~prog_clock_reg[0];
	end

// ----- End raw programming clock signal generation -----

// ----- Actual programming clock is triggered only when config_done and prog_reset are disabled -----
	assign prog_clock[0] = prog_clock_reg[0] & (~config_done[0]) & (~prog_reset[0]);

// ----- Begin raw operating clock signal generation -----
initial
	begin
		op_clock_reg[0] = {1{1'b0}};
	end
always wait(~greset)
	begin
		#0.558185935	op_clock_reg[0] = ~op_clock_reg[0];
	end

// ----- End raw operating clock signal generation -----
// ----- Actual operating clock is triggered only when config_done is enabled -----
	assign op_clock[0] = op_clock_reg[0] & config_done[0];

// ----- Begin programming reset signal generation -----
initial
	begin
		prog_reset[0] = {1{1'b1}};
	#10	prog_reset[0] = {1{1'b0}};
	end

// ----- End programming reset signal generation -----

// ----- Begin programming set signal generation: always disabled -----
initial
	begin
		prog_set[0] = {1{1'b0}};
	end

// ----- End programming set signal generation: always disabled -----

// ----- Begin operating reset signal generation -----
// ----- Reset signal is enabled until the first clock cycle in operation phase -----
initial
	begin
		greset[0] = {1{1'b1}};
	wait(config_done)
	#1.11637187	greset[0] = {1{1'b1}};
	#2.23274374	greset[0] = {1{1'b0}};
	end

// ----- End operating reset signal generation -----
// ----- Begin operating set signal generation: always disabled -----
initial
	begin
		gset[0] = {1{1'b0}};
	end

// ----- End operating set signal generation: always disabled -----

// ----- Begin connecting global ports of FPGA fabric to stimuli -----
	assign clk[0] = op_clock[0];
	assign prog_clk[0] = prog_clock[0];
	assign reset[0] = greset[0];
	assign pReset[0] = prog_reset[0];
	assign set[0] = gset[0];
// ----- End connecting global ports of FPGA fabric to stimuli -----
// ----- FPGA top-level module to be capsulated -----
	fpga_top FPGA_DUT (
		.pReset(pReset[0]),
		.prog_clk(prog_clk[0]),
		.set(set[0]),
		.reset(reset[0]),
		.clk(clk[0]),
		.gfpga_pad_iopad_pad(gfpga_pad_iopad_pad[0:63]),
		.ccff_head(ccff_head[0]),
		.ccff_tail(ccff_tail[0]));

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input a is mapped to FPGA IOPAD gfpga_pad_iopad_pad[17] -----
	assign gfpga_pad_iopad_pad[17] = a[0];
// ----- Blif Benchmark input b is mapped to FPGA IOPAD gfpga_pad_iopad_pad[40] -----
	assign gfpga_pad_iopad_pad[40] = b[0];
// ----- Blif Benchmark output out_c is mapped to FPGA IOPAD gfpga_pad_iopad_pad[46] -----
	assign out_c_fpga[0] = gfpga_pad_iopad_pad[46];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_iopad_pad[0] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[1] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[2] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[3] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[4] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[5] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[6] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[7] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[8] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[9] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[10] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[11] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[12] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[13] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[14] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[15] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[16] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[18] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[19] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[20] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[21] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[22] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[23] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[24] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[25] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[26] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[27] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[28] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[29] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[30] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[31] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[32] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[33] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[34] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[35] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[36] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[37] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[38] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[39] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[41] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[42] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[43] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[44] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[45] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[47] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[48] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[49] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[50] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[51] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[52] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[53] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[54] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[55] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[56] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[57] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[58] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[59] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[60] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[61] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[62] = {1{1'b0}};
	assign gfpga_pad_iopad_pad[63] = {1{1'b0}};

`ifdef AUTOCHECKED_SIMULATION
// ----- Reference Benchmark Instanication -------
	and2 REF_DUT(
		.a(a),
		.b(b),
		.c(out_c_benchmark)	);
// ----- End reference Benchmark Instanication -------

`endif


// ----- Task: input values during a programming clock cycle -----
task prog_cycle_task;
input [0:0] ccff_head_val;
	begin
		@(negedge prog_clock[0]);
			ccff_head[0] = ccff_head_val[0];
	end
endtask

// ----- Begin bitstream loading during configuration phase -----
initial
	begin
// ----- Configuration chain default input -----
		ccff_head[0] = {1{1'b0}};
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		@(negedge prog_clock[0]);
			config_done[0] <= {1{1'b1}};
	end
// ----- End bitstream loading during configuration phase -----
// ----- Input Initialization -------
	initial begin
		a <= 1'b0;
		b <= 1'b0;

		out_c_flag[0] <= 1'b0;
	end

// ----- Input Stimulus -------
	always@(negedge op_clock[0]) begin
		a <= $random;
		b <= $random;
	end

`ifdef AUTOCHECKED_SIMULATION
// ----- Begin checking output vectors -------
// ----- Skip the first falling edge of clock, it is for initialization -------
	reg [0:0] sim_start;

	always@(negedge op_clock[0]) begin
		if (1'b1 == sim_start[0]) begin
			sim_start[0] <= ~sim_start[0];
		end else begin
			if(!(out_c_fpga === out_c_benchmark) && !(out_c_benchmark === 1'bx)) begin
				out_c_flag <= 1'b1;
			end else begin
				out_c_flag<= 1'b0;
			end
		end
	end

	always@(posedge out_c_flag) begin
		if(out_c_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out_c_fpga at time = %t", $realtime);
		end
	end

`endif

`ifdef ICARUS_SIMULATOR
// ----- Begin Icarus requirement -------
	initial begin
		$dumpfile("and2_formal.vcd");
		$dumpvars(1, and2_autocheck_top_tb);
	end
`endif
// ----- END Icarus requirement -------

initial begin
	sim_start[0] <= 1'b1;
	$timeformat(-9, 2, "ns", 20);
	$display("Simulation start");
// ----- Can be changed by the user for his/her need -------
	#18792
	if(nb_error == 0) begin
		$display("Simulation Succeed");
	end else begin
		$display("Simulation Failed with %d error(s)", nb_error);
	end
	$finish;
end

endmodule
// ----- END Verilog module for and2_autocheck_top_tb -----

